package pmd901_bus_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "pmd901_bus_trans.sv"
`include "pmd901_bus_agent_config.sv"

`include "pmd901_bus_monitor.sv"
`include "pmd901_bus_driver.sv"
`include "pmd901_bus_sequencer.sv"

`include "pmd901_bus_recorder.sv"

`include "pmd901_bus_agent.sv"

// API sequences
`include "pmd901_sequences/pmd901_bus_enable_sequence.sv"
`include "pmd901_sequences/pmd901_bus_bending_sequence.sv"
`include "pmd901_sequences/pmd901_bus_speed_sequence.sv"
`include "pmd901_sequences/pmd901_bus_rand_speed_bending_sequence.sv"
endpackage 
