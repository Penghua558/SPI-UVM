package pmd901_bus_sequence_lib_pkg;
    `include "./pmd901_sequences/pmd901_bus_enable_sequence.sv"
    `include "./pmd901_sequences/pmd901_bus_bending_sequence.sv"
    `include "./pmd901_sequences/pmd901_bus_speed_sequence.sv"
endpackage: pmd901_bus_sequence_lib_pkg
