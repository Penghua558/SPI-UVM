package testcase_lib_pkg;

// Standard UVM import & include:
import uvm_pkg::*;
`include "uvm_macros.svh"

import env_pkg::*;
import pmd901_agent_pkg::*;
import apb_agent_pkg::*;
import spi_bus_sequence_lib_pkg::*;
import spi_reg_pkg::*;

// testcases
`include "test_base.sv"
`include "test.sv"

endpackage: testcase_lib_pkg
