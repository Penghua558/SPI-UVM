package pmd901_bus_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "pmd901_bus_trans.sv"
`include "pmd901_bus_agent_config.sv"

`include "pmd901_bus_driver.sv"
`include "pmd901_bus_sequencer.sv"
`include "pmd901_bus_sequence.sv"

`include "pmd901_bus_agent.sv"
endpackage 
