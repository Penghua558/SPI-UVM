package pmd901_bus_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "pmd901_bus_trans.sv"
`include "pmd901_bus_agent_config.sv"

`include "pmd901_bus_monitor.sv"
`include "pmd901_bus_driver.sv"
`include "pmd901_bus_sequencer.sv"

import pmd901_bus_sequence_lib_pkg::*;

`include "pmd901_bus_agent.sv"
endpackage 
