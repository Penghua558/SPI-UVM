import apb_agent_dec::*;
class apb_rand_read_sequence extends uvm_sequence #(apb_trans);

// UVM Factory Registration Macro
//
`uvm_object_utils(apb_rand_read_sequence)


//------------------------------------------
// Data Members (Outputs rand, inputs non-rand)
//------------------------------------------
logic [15:0] data;

//------------------------------------------
// Constraints
//------------------------------------------



//------------------------------------------
// Methods
//------------------------------------------

// Standard UVM Methods:
extern function new(string name = "apb_rand_read_sequence");
extern task body;
extern task read(uvm_sequencer_base seqr, uvm_sequencer_base parent = null);

endclass:apb_rand_read_sequence

function apb_rand_read_sequence::new(string name = "apb_rand_read_sequence");
  super.new(name);
endfunction

task apb_rand_read_sequence::body;
    apb_agent_config m_cfg = apb_agent_config::get_config(this);
    apb_trans req = apb_trans::type_id::create("req");;

    begin
        start_item(req);
        assert(req.randomize() with {
            wr == READ;
            addr >= m_cfg.start_address[m_cfg.apb_index]; 
            addr <= m_cfg.start_address[m_cfg.apb_index] + 
                m_cfg.range[m_cfg.apb_index];
        });
        finish_item(req);
        data = req.rdata;
    end
endtask:body

task apb_rand_read_sequence::read(uvm_sequencer_base seqr, 
    uvm_sequencer_base parent = null);
    this.start(seqr, parent);
endtask
