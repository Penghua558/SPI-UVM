package pmd901_bus_sequence_lib_pkg;
endpackage: pmd901_bus_sequence_lib_pkg
