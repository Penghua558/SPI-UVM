package pmd901_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "pmd901_trans.sv"
`include "pmd901_agent_config.sv"

`include "pmd901_monitor.sv"
`include "pmd901_driver.sv"
`include "pmd901_sequencer.sv"
`include "pmd901_sequence.sv"

`include "pmd901_agent.sv"
endpackage: pmd901_agent_pkg 
