//
//------------------------------------------------------------------------------
//   Copyright 2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------
//
//------------------------------------------------------------------------------
//   Copyright 2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------
//----------------------------------------------------------------------
//   THIS IS AUTOMATICALLY GENERATED CODE
//   Generated by Mentor Graphics' Register Assistant UVM V4.6 (Build 8)
//   UVM Register Kit version 1.1
//----------------------------------------------------------------------
// Project         : register_model
// Unit            : spi_reg_pkg
// File            : spi_reg_pkg.sv
//----------------------------------------------------------------------
// Created by      : cgales
// Creation Date   : 2/19/16 3:24 PM
//----------------------------------------------------------------------
// Title           : register_model
//
// Description     : 
//
//----------------------------------------------------------------------

//----------------------------------------------------------------------
// spi_reg_pkg
//----------------------------------------------------------------------
package spi_reg_pkg;

   import uvm_pkg::*;

   `include "uvm_macros.svh"

   /* DEFINE REGISTER CLASSES */



   //--------------------------------------------------------------------
   // Class: divider_reg
   // 
   // Divider
   //--------------------------------------------------------------------

   class divider_reg extends uvm_reg;
      `uvm_object_utils(divider_reg)

      rand uvm_reg_field ratio; 


      // Function: coverage
      // 
      covergroup cg_vals;
         ratio	 : coverpoint ratio.value[15:0];
      endgroup



      // Function: new
      // 
      function new(string name = "divider_reg");
         super.new(name, 32, build_coverage(UVM_CVR_FIELD_VALS));
         add_coverage(build_coverage(UVM_CVR_FIELD_VALS));
         if(has_coverage(UVM_CVR_FIELD_VALS))
            cg_vals = new();
      endfunction


      // Function: sample_values
      // 
      virtual function void sample_values();
         super.sample_values();
         if (get_coverage(UVM_CVR_FIELD_VALS))
            cg_vals.sample();
      endfunction


      // Function: build
      // 
      virtual function void build();
         ratio = uvm_reg_field::type_id::create("ratio");

         ratio.configure(this, 16, 0, "RW", 0, 16'h0000, 1, 1, 1);
      endfunction
   endclass



   //--------------------------------------------------------------------
   // Class: rxtx0_reg
   // 
   // RXTX0
   //--------------------------------------------------------------------

   class rxtx0_reg extends uvm_reg;
      `uvm_object_utils(rxtx0_reg)

      rand uvm_reg_field F;


      // Function: new
      // 
      function new(string name = "rxtx0_reg");
         super.new(name, 32, UVM_NO_COVERAGE);
      endfunction


      // Function: build
      // 
      virtual function void build();
         F = uvm_reg_field::type_id::create("F");
         F.configure(this, 32, 0, "RW", 1, 32'h00000000, 1, 1, 1);
      endfunction
   endclass



   //--------------------------------------------------------------------
   // Class: rxtx3_reg
   // 
   // RXTX3
   //--------------------------------------------------------------------

   class rxtx3_reg extends uvm_reg;
      `uvm_object_utils(rxtx3_reg)

      rand uvm_reg_field F;


      // Function: new
      // 
      function new(string name = "rxtx3_reg");
         super.new(name, 32, UVM_NO_COVERAGE);
      endfunction


      // Function: build
      // 
      virtual function void build();
         F = uvm_reg_field::type_id::create("F");
         F.configure(this, 32, 0, "RW", 1, 32'h00000000, 1, 1, 1);
      endfunction
   endclass



   //--------------------------------------------------------------------
   // Class: rxtx1_reg
   // 
   // RXTX1
   //--------------------------------------------------------------------

   class rxtx1_reg extends uvm_reg;
      `uvm_object_utils(rxtx1_reg)

      rand uvm_reg_field F;


      // Function: new
      // 
      function new(string name = "rxtx1_reg");
         super.new(name, 32, UVM_NO_COVERAGE);
      endfunction


      // Function: build
      // 
      virtual function void build();
         F = uvm_reg_field::type_id::create("F");
         F.configure(this, 32, 0, "RW", 1, 32'h00000000, 1, 1, 1);
      endfunction
   endclass



   //--------------------------------------------------------------------
   // Class: ss_reg
   // 
   // Status
   //--------------------------------------------------------------------

   class ss_reg extends uvm_reg;
      `uvm_object_utils(ss_reg)

      rand uvm_reg_field reserved; 
      rand uvm_reg_field cs; 


      // Function: coverage
      // 
      covergroup cg_vals;
         cs	 : coverpoint cs.value[7:0];
      endgroup



      // Function: new
      // 
      function new(string name = "ss_reg");
         super.new(name, 32, build_coverage(UVM_CVR_FIELD_VALS));
         add_coverage(build_coverage(UVM_CVR_FIELD_VALS));
         if(has_coverage(UVM_CVR_FIELD_VALS))
            cg_vals = new();
      endfunction


      // Function: sample_values
      // 
      virtual function void sample_values();
         super.sample_values();
         if (get_coverage(UVM_CVR_FIELD_VALS))
            cg_vals.sample();
      endfunction


      // Function: build
      // 
      virtual function void build();
         reserved = uvm_reg_field::type_id::create("reserved");
         cs = uvm_reg_field::type_id::create("cs");

         reserved.configure(this, 8, 8, "RW", 0, 8'h00, 1, 1, 1);
         cs.configure(this, 8, 0, "RW", 0, 8'h00, 1, 1, 1);
      endfunction
   endclass



   //--------------------------------------------------------------------
   // Class: rxtx2_reg
   // 
   // RXTX2
   //--------------------------------------------------------------------

   class rxtx2_reg extends uvm_reg;
      `uvm_object_utils(rxtx2_reg)

      rand uvm_reg_field F;


      // Function: new
      // 
      function new(string name = "rxtx2_reg");
         super.new(name, 32, UVM_NO_COVERAGE);
      endfunction


      // Function: build
      // 
      virtual function void build();
         F = uvm_reg_field::type_id::create("F");
         F.configure(this, 32, 0, "RW", 1, 32'h00000000, 1, 1, 1);
      endfunction
   endclass



   //--------------------------------------------------------------------
   // Class: ctrl_reg
   // 
   // Control Status Register
   //--------------------------------------------------------------------

   class ctrl_reg extends uvm_reg;
      `uvm_object_utils(ctrl_reg)

      rand uvm_reg_field ass; 
      rand uvm_reg_field ie; 
      rand uvm_reg_field lsb; 
      rand uvm_reg_field tx_neg; 
      rand uvm_reg_field rx_neg; 
      rand uvm_reg_field go_bsy; 
      rand uvm_reg_field reserved2; 
      rand uvm_reg_field char_len; 


      // Function: coverage
      // 
      covergroup cg_vals;
         ass	 : coverpoint ass.value[0];
         ie	 : coverpoint ie.value[0];
         lsb	 : coverpoint lsb.value[0];
         tx_neg	 : coverpoint tx_neg.value[0];
         rx_neg	 : coverpoint rx_neg.value[0];
         go_bsy	 : coverpoint go_bsy.value[0];
         char_len	 : coverpoint char_len.value[6:0];
      endgroup



      // Function: new
      // 
      function new(string name = "ctrl_reg");
         super.new(name, 32, build_coverage(UVM_CVR_FIELD_VALS));
         add_coverage(build_coverage(UVM_CVR_FIELD_VALS));
         if(has_coverage(UVM_CVR_FIELD_VALS))
            cg_vals = new();
      endfunction


      // Function: sample_values
      // 
      virtual function void sample_values();
         super.sample_values();
         if (get_coverage(UVM_CVR_FIELD_VALS))
            cg_vals.sample();
      endfunction


      // Function: build
      // 
      virtual function void build();
         ass = uvm_reg_field::type_id::create("ass");
         ie = uvm_reg_field::type_id::create("ie");
         lsb = uvm_reg_field::type_id::create("lsb");
         tx_neg = uvm_reg_field::type_id::create("tx_neg");
         rx_neg = uvm_reg_field::type_id::create("rx_neg");
         go_bsy = uvm_reg_field::type_id::create("go_bsy");
         reserved2 = uvm_reg_field::type_id::create("reserved2");
         char_len = uvm_reg_field::type_id::create("char_len");

         ass.configure(this, 1, 13, "RW", 0, 1'b0, 1, 1, 0);
         ie.configure(this, 1, 12, "RW", 0, 1'b0, 1, 1, 0);
         lsb.configure(this, 1, 11, "RW", 0, 1'b0, 1, 1, 0);
         tx_neg.configure(this, 1, 10, "RW", 0, 1'b0, 1, 1, 0);
         rx_neg.configure(this, 1, 9, "RW", 0, 1'b0, 1, 1, 0);
         go_bsy.configure(this, 1, 8, "RW", 0, 1'b0, 1, 1, 0);
         reserved2.configure(this, 1, 7, "RW", 0, 1'b0, 1, 1, 0);
         char_len.configure(this, 7, 0, "RW", 0, 7'b0000000, 1, 1, 0);
      endfunction
   endclass




   /* BLOCKS */



   //--------------------------------------------------------------------
   // Class: spi_reg_block
   // 
   //--------------------------------------------------------------------

   class spi_reg_block extends uvm_reg_block;
      `uvm_object_utils(spi_reg_block)

      rand rxtx0_reg rxtx0; // RXTX0
      rand rxtx1_reg rxtx1; // RXTX1
      rand rxtx2_reg rxtx2; // RXTX2
      rand rxtx3_reg rxtx3; // RXTX3
      rand ctrl_reg ctrl; // Control Status Register
      rand divider_reg divider; // Divider
      rand ss_reg ss; // Status

      uvm_reg_map spi_reg_block_map; 


      // Function: new
      // 
      function new(string name = "spi_reg_block");
         super.new(name, build_coverage(UVM_CVR_ALL));
      endfunction


      // Function: build
      // 
      virtual function void build();
         rxtx0 = rxtx0_reg::type_id::create("rxtx0");
         rxtx0.configure(this);
         rxtx0.build();

         rxtx1 = rxtx1_reg::type_id::create("rxtx1");
         rxtx1.configure(this);
         rxtx1.build();

         rxtx2 = rxtx2_reg::type_id::create("rxtx2");
         rxtx2.configure(this);
         rxtx2.build();

         rxtx3 = rxtx3_reg::type_id::create("rxtx3");
         rxtx3.configure(this);
         rxtx3.build();

         ctrl = ctrl_reg::type_id::create("ctrl");
         ctrl.configure(this);
         ctrl.build();

         divider = divider_reg::type_id::create("divider");
         divider.configure(this);
         divider.build();

         ss = ss_reg::type_id::create("ss");
         ss.configure(this);
         ss.build();

         spi_reg_block_map = create_map("spi_reg_block_map", 'h0, 4, UVM_LITTLE_ENDIAN, 1);
         default_map = spi_reg_block_map;

         spi_reg_block_map.add_reg(rxtx0, 'h0, "RW");
         spi_reg_block_map.add_reg(rxtx1, 'h4, "RW");
         spi_reg_block_map.add_reg(rxtx2, 'h8, "RW");
         spi_reg_block_map.add_reg(rxtx3, 'hc, "RW");
         spi_reg_block_map.add_reg(ctrl, 'h10, "RW");
         spi_reg_block_map.add_reg(divider, 'h14, "RW");
         spi_reg_block_map.add_reg(ss, 'h18, "RW");

         lock_model();
      endfunction
   endclass


endpackage
