package pmd901_agent_dec;
    typedef enum {
        POWER_DOWN,
        NORMAL_WORKING,
        BENDING_WORKING
        } work_status_e;
endpackage: pmd901_agent_dec
